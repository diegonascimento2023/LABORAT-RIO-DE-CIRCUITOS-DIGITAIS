module seteSeg (s, hex);
	input [3:0] s;
	output [6:0] hex;

	assign hex =(s == 4'b0000)? 7'b100_0000:	// 0
					(s == 4'b0001)? 7'b111_1001:	// 1
					(s == 4'b0010)? 7'b010_0100:	// 2
					(s == 4'b0011)? 7'b011_0000:	// 3
					(s == 4'b0100)? 7'b001_1001:	// 4
					(s == 4'b0101)? 7'b001_0010:	// 5
					(s == 4'b0110)? 7'b000_0010:	// 6
					(s == 4'b0111)? 7'b111_1000:	// 7
					(s == 4'b1000)? 7'b000_0000:	// 8
					(s == 4'b1001)? 7'b001_1000:	// 9
					7'b111_1111; // Null
endmodule
